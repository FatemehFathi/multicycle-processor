`timescale 1ns/1ns

module AND(input a, b, output w);
  assign w = a & b;
endmodule




module OR(input a, b, output w);
  assign w = a | b;
endmodule

